library verilog;
use verilog.vl_types.all;
entity test_sequences_define_sv_unit is
end test_sequences_define_sv_unit;
