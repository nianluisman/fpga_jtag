// Define IDCODE Value
`define IDCODE_VALUE  32'h149511c3

// Length of the Instruction register
`define	IR_LENGTH	4

`define IDCODE          4'b0010